library verilog;
use verilog.vl_types.all;
entity bitdetector_tb is
end bitdetector_tb;
