library verilog;
use verilog.vl_types.all;
entity testbit is
end testbit;
